library ieee;
use ieee.std_logic_1164.all;

entity neorv32_cfs is
    generic (
        CFS_CONFIG : std_ulogic_vector(31 downto 0);
        CFS_IN_SIZE : natural;
        CFS_OUT_SIZE : natural
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        bus_req_i : in bus_req_t;
        bus_rsp_o : out bus_rsp_t;
        clkgen_en_o : out std_ulogic;
        clkgen_i : in std_ulogic_vector(7 downto 0);
        irq_o : out std_ulogic;
        cfs_in_i : in std_ulogic_vector(CFS_IN_SIZE-1 downto 0);
        cfs_out_o : out std_ulogic_vector(CFS_OUT_SIZE-1 downto 0)
    );
end entity neorv32_cfs;