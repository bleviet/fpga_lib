library ieee;
use ieee.std_logic_1164.all;

entity neorv32_uart is
    generic (
        SIM_MODE_EN : boolean;
        SIM_LOG_FILE : string;
        UART_RX_FIFO : natural range 1 to 2**15;
        UART_TX_FIFO : natural range 1 to 2**15
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        bus_req_i : in bus_req_t;
        bus_rsp_o : out bus_rsp_t;
        clkgen_en_o : out std_ulogic;
        clkgen_i : in std_ulogic_vector(7 downto 0);
        uart_txd_o : out std_ulogic;
        uart_rxd_i : in std_ulogic;
        uart_rtsn_o : out std_ulogic;
        uart_ctsn_i : in std_ulogic;
        irq_rx_o : out std_ulogic;
        irq_tx_o : out std_ulogic
    );
end entity neorv32_uart;