library ieee;
use ieee.std_logic_1164.all;

entity neorv32_top is
    generic (
        CLOCK_FREQUENCY : natural := 0;
        HART_BASE : natural := 0;
        DUAL_CORE_EN : boolean := false;
        BOOT_MODE_SELECT : natural range 0 to 2 := 0;
        BOOT_ADDR_CUSTOM : std_ulogic_vector(31 downto 0) := x"00000000";
        OCD_EN : boolean := false;
        OCD_HW_BREAKPOINT : boolean := false;
        OCD_AUTHENTICATION : boolean := false;
        OCD_JEDEC_ID : std_ulogic_vector(10 downto 0) := "00000000000";
        RISCV_ISA_C : boolean := false;
        RISCV_ISA_E : boolean := false;
        RISCV_ISA_M : boolean := false;
        RISCV_ISA_U : boolean := false;
        RISCV_ISA_Zaamo : boolean := false;
        RISCV_ISA_Zalrsc : boolean := false;
        RISCV_ISA_Zba : boolean := false;
        RISCV_ISA_Zbb : boolean := false;
        RISCV_ISA_Zbkb : boolean := false;
        RISCV_ISA_Zbkc : boolean := false;
        RISCV_ISA_Zbkx : boolean := false;
        RISCV_ISA_Zbs : boolean := false;
        RISCV_ISA_Zfinx : boolean := false;
        RISCV_ISA_Zicntr : boolean := false;
        RISCV_ISA_Zicond : boolean := false;
        RISCV_ISA_Zihpm : boolean := false;
        RISCV_ISA_Zknd : boolean := false;
        RISCV_ISA_Zkne : boolean := false;
        RISCV_ISA_Zknh : boolean := false;
        RISCV_ISA_Zksed : boolean := false;
        RISCV_ISA_Zksh : boolean := false;
        RISCV_ISA_Zmmul : boolean := false;
        RISCV_ISA_Zxcfu : boolean := false;
        CPU_FAST_MUL_EN : boolean := false;
        CPU_FAST_SHIFT_EN : boolean := false;
        CPU_RF_HW_RST_EN : boolean := false;
        PMP_NUM_REGIONS : natural range 0 to 16 := 0;
        PMP_MIN_GRANULARITY : natural := 4;
        PMP_TOR_MODE_EN : boolean := false;
        PMP_NAP_MODE_EN : boolean := false;
        HPM_NUM_CNTS : natural range 0 to 13 := 0;
        HPM_CNT_WIDTH : natural range 0 to 64 := 40;
        MEM_INT_IMEM_EN : boolean := false;
        MEM_INT_IMEM_SIZE : natural := 16*1024;
        MEM_INT_DMEM_EN : boolean := false;
        MEM_INT_DMEM_SIZE : natural := 8*1024;
        ICACHE_EN : boolean := false;
        ICACHE_NUM_BLOCKS : natural range 1 to 256 := 4;
        ICACHE_BLOCK_SIZE : natural range 4 to 2**16 := 64;
        DCACHE_EN : boolean := false;
        DCACHE_NUM_BLOCKS : natural range 1 to 256 := 4;
        DCACHE_BLOCK_SIZE : natural range 4 to 2**16 := 64;
        XBUS_EN : boolean := false;
        XBUS_TIMEOUT : natural := 255;
        XBUS_REGSTAGE_EN : boolean := false;
        XBUS_CACHE_EN : boolean := false;
        XBUS_CACHE_NUM_BLOCKS : natural range 1 to 256 := 64;
        XBUS_CACHE_BLOCK_SIZE : natural range 1 to 2**16 := 32;
        IO_DISABLE_SYSINFO : boolean := false;
        IO_GPIO_NUM : natural range 0 to 32 := 0;
        IO_CLINT_EN : boolean := false;
        IO_UART0_EN : boolean := false;
        IO_UART0_RX_FIFO : natural range 1 to 2**15 := 1;
        IO_UART0_TX_FIFO : natural range 1 to 2**15 := 1;
        IO_UART1_EN : boolean := false;
        IO_UART1_RX_FIFO : natural range 1 to 2**15 := 1;
        IO_UART1_TX_FIFO : natural range 1 to 2**15 := 1;
        IO_SPI_EN : boolean := false;
        IO_SPI_FIFO : natural range 1 to 2**15 := 1;
        IO_SDI_EN : boolean := false;
        IO_SDI_FIFO : natural range 1 to 2**15 := 1;
        IO_TWI_EN : boolean := false;
        IO_TWI_FIFO : natural range 1 to 2**15 := 1;
        IO_TWD_EN : boolean := false;
        IO_TWD_RX_FIFO : natural range 1 to 2**15 := 1;
        IO_TWD_TX_FIFO : natural range 1 to 2**15 := 1;
        IO_PWM_NUM_CH : natural range 0 to 16 := 0;
        IO_WDT_EN : boolean := false;
        IO_TRNG_EN : boolean := false;
        IO_TRNG_FIFO : natural range 1 to 2**15 := 1;
        IO_CFS_EN : boolean := false;
        IO_CFS_CONFIG : std_ulogic_vector(31 downto 0) := x"00000000";
        IO_CFS_IN_SIZE : natural := 32;
        IO_CFS_OUT_SIZE : natural := 32;
        IO_NEOLED_EN : boolean := false;
        IO_NEOLED_TX_FIFO : natural range 1 to 2**15 := 1;
        IO_GPTMR_EN : boolean := false;
        IO_ONEWIRE_EN : boolean := false;
        IO_ONEWIRE_FIFO : natural range 1 to 2**15 := 1;
        IO_DMA_EN : boolean := false;
        IO_SLINK_EN : boolean := false;
        IO_SLINK_RX_FIFO : natural range 1 to 2**15 := 1;
        IO_SLINK_TX_FIFO : natural range 1 to 2**15 := 1;
        IO_CRC_EN : boolean := false;
        IO_HWSPINLOCK_EN : boolean := false
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        rstn_ocd_o : out std_ulogic;
        rstn_wdt_o : out std_ulogic;
        jtag_tck_i : in std_ulogic := 'L';
        jtag_tdi_i : in std_ulogic := 'L';
        jtag_tdo_o : out std_ulogic;
        jtag_tms_i : in std_ulogic := 'L';
        xbus_adr_o : out std_ulogic_vector(31 downto 0);
        xbus_dat_o : out std_ulogic_vector(31 downto 0);
        xbus_tag_o : out std_ulogic_vector(2 downto 0);
        xbus_we_o : out std_ulogic;
        xbus_sel_o : out std_ulogic_vector(3 downto 0);
        xbus_stb_o : out std_ulogic;
        xbus_cyc_o : out std_ulogic;
        xbus_dat_i : in std_ulogic_vector(31 downto 0) := (others => 'L');
        xbus_ack_i : in std_ulogic := 'L';
        xbus_err_i : in std_ulogic := 'L';
        slink_rx_dat_i : in std_ulogic_vector(31 downto 0) := (others => 'L');
        slink_rx_src_i : in std_ulogic_vector(3 downto 0)  := (others => 'L');
        slink_rx_val_i : in std_ulogic := 'L';
        slink_rx_lst_i : in std_ulogic := 'L';
        slink_rx_rdy_o : out std_ulogic;
        slink_tx_dat_o : out std_ulogic_vector(31 downto 0);
        slink_tx_dst_o : out std_ulogic_vector(3 downto 0);
        slink_tx_val_o : out std_ulogic;
        slink_tx_lst_o : out std_ulogic;
        slink_tx_rdy_i : in std_ulogic := 'L';
        gpio_o : out std_ulogic_vector(31 downto 0);
        gpio_i : in std_ulogic_vector(31 downto 0) := (others => 'L');
        uart0_txd_o : out std_ulogic;
        uart0_rxd_i : in std_ulogic := 'L';
        uart0_rtsn_o : out std_ulogic;
        uart0_ctsn_i : in std_ulogic := 'L';
        uart1_txd_o : out std_ulogic;
        uart1_rxd_i : in std_ulogic := 'L';
        uart1_rtsn_o : out std_ulogic;
        uart1_ctsn_i : in std_ulogic := 'L';
        spi_clk_o : out std_ulogic;
        spi_dat_o : out std_ulogic;
        spi_dat_i : in std_ulogic := 'L';
        spi_csn_o : out std_ulogic_vector(7 downto 0);
        sdi_clk_i : in std_ulogic := 'L';
        sdi_dat_o : out std_ulogic;
        sdi_dat_i : in std_ulogic := 'L';
        sdi_csn_i : in std_ulogic := 'H';
        twi_sda_i : in std_ulogic := 'H';
        twi_sda_o : out std_ulogic;
        twi_scl_i : in std_ulogic := 'H';
        twi_scl_o : out std_ulogic;
        twd_sda_i : in std_ulogic := 'H';
        twd_sda_o : out std_ulogic;
        twd_scl_i : in std_ulogic := 'H';
        twd_scl_o : out std_ulogic;
        onewire_i : in std_ulogic := 'H';
        onewire_o : out std_ulogic;
        pwm_o : out std_ulogic_vector(15 downto 0);
        cfs_in_i : in std_ulogic_vector(IO_CFS_IN_SIZE-1 downto 0) := (others => 'L');
        cfs_out_o : out std_ulogic_vector(IO_CFS_OUT_SIZE-1 downto 0);
        neoled_o : out std_ulogic;
        mtime_time_o : out std_ulogic_vector(63 downto 0);
        mtime_irq_i : in std_ulogic := 'L';
        msw_irq_i : in std_ulogic := 'L';
        mext_irq_i : in std_ulogic := 'L'
    );
end entity neorv32_top;