library ieee;
use ieee.std_logic_1164.all;

entity neorv32_cpu_alu is
    generic (
        RISCV_ISA_M : boolean;
        RISCV_ISA_Zba : boolean;
        RISCV_ISA_Zbb : boolean;
        RISCV_ISA_Zbkb : boolean;
        RISCV_ISA_Zbkc : boolean;
        RISCV_ISA_Zbkx : boolean;
        RISCV_ISA_Zbs : boolean;
        RISCV_ISA_Zfinx : boolean;
        RISCV_ISA_Zicond : boolean;
        RISCV_ISA_Zknd : boolean;
        RISCV_ISA_Zkne : boolean;
        RISCV_ISA_Zknh : boolean;
        RISCV_ISA_Zksed : boolean;
        RISCV_ISA_Zksh : boolean;
        RISCV_ISA_Zmmul : boolean;
        RISCV_ISA_Zxcfu : boolean;
        FAST_MUL_EN : boolean;
        FAST_SHIFT_EN : boolean
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        ctrl_i : in ctrl_bus_t;
        rs1_i : in std_ulogic_vector(XLEN-1 downto 0);
        rs2_i : in std_ulogic_vector(XLEN-1 downto 0);
        rs3_i : in std_ulogic_vector(XLEN-1 downto 0);
        cmp_o : out std_ulogic_vector(1 downto 0);
        res_o : out std_ulogic_vector(XLEN-1 downto 0);
        add_o : out std_ulogic_vector(XLEN-1 downto 0);
        csr_o : out std_ulogic_vector(XLEN-1 downto 0);
        done_o : out std_ulogic
    );
end entity neorv32_cpu_alu;