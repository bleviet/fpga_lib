library ieee;
use ieee.std_logic_1164.all;

entity neorv32_cpu_lsu is
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic := '0';
        ctrl_i : in ctrl_bus_t;
        addr_i : in std_ulogic_vector(XLEN-1 downto 0);
        wdata_i : in std_ulogic_vector(XLEN-1 downto 0);
        rdata_o : out std_ulogic_vector(XLEN-1 downto 0);
        mar_o : out std_ulogic_vector(XLEN-1 downto 0);
        wait_o : out std_ulogic;
        err_o : out std_ulogic_vector(3 downto 0);
        pmp_fault_i : in std_ulogic;
        dbus_req_o : out bus_req_t;
        dbus_rsp_i : in bus_rsp_t
    );
end entity neorv32_cpu_lsu;