library ieee;
use ieee.std_logic_1164.all;

entity neorv32_xbus is
    generic (
        TIMEOUT_VAL : natural;
        REGSTAGE_EN : boolean
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        bus_req_i : in bus_req_t;
        bus_rsp_o : out bus_rsp_t;
        xbus_adr_o : out std_ulogic_vector(31 downto 0);
        xbus_dat_i : in std_ulogic_vector(31 downto 0);
        xbus_dat_o : out std_ulogic_vector(31 downto 0);
        xbus_tag_o : out std_ulogic_vector(2 downto 0);
        xbus_we_o : out std_ulogic;
        xbus_sel_o : out std_ulogic_vector(3 downto 0);
        xbus_stb_o : out std_ulogic;
        xbus_cyc_o : out std_ulogic;
        xbus_ack_i : in std_ulogic;
        xbus_err_i : in std_ulogic
    );
end entity neorv32_xbus;