library ieee;
use ieee.std_logic_1164.all;

entity neorv32_cpu_cp_bitmanip is
    generic (
        EN_FAST_SHIFT : boolean;
        EN_ZBA : boolean;
        EN_ZBB : boolean;
        EN_ZBKC : boolean;
        EN_ZBKB : boolean;
        EN_ZBS : boolean
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        ctrl_i : in ctrl_bus_t;
        cmp_i : in std_ulogic_vector(1 downto 0);
        rs1_i : in std_ulogic_vector(XLEN-1 downto 0);
        rs2_i : in std_ulogic_vector(XLEN-1 downto 0);
        shamt_i : in std_ulogic_vector(index_size_f(XLEN)-1 downto 0);
        res_o : out std_ulogic_vector(XLEN-1 downto 0);
        valid_o : out std_ulogic
    );
end entity neorv32_cpu_cp_bitmanip;