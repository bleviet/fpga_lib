library ieee;
use ieee.std_logic_1164.all;

entity neorv32_bus_switch is
    generic (
        ROUND_ROBIN_EN : boolean := false;
        PORT_A_READ_ONLY : boolean := false;
        PORT_B_READ_ONLY : boolean := false
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        a_req_i : in bus_req_t;
        a_rsp_o : out bus_rsp_t;
        b_req_i : in bus_req_t;
        b_rsp_o : out bus_rsp_t;
        x_req_o : out bus_req_t;
        x_rsp_i : in bus_rsp_t
    );
end entity neorv32_bus_switch;