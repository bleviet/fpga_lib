library ieee;
use ieee.std_logic_1164.all;

entity neorv32_cpu_control is
    generic (
        HART_ID : natural range 0 to 1023;
        BOOT_ADDR : std_ulogic_vector(31 downto 0);
        DEBUG_PARK_ADDR : std_ulogic_vector(31 downto 0);
        DEBUG_EXC_ADDR : std_ulogic_vector(31 downto 0);
        RISCV_ISA_A : boolean;
        RISCV_ISA_B : boolean;
        RISCV_ISA_C : boolean;
        RISCV_ISA_E : boolean;
        RISCV_ISA_M : boolean;
        RISCV_ISA_U : boolean;
        RISCV_ISA_Zaamo : boolean;
        RISCV_ISA_Zalrsc : boolean;
        RISCV_ISA_Zba : boolean;
        RISCV_ISA_Zbb : boolean;
        RISCV_ISA_Zbkb : boolean;
        RISCV_ISA_Zbkc : boolean;
        RISCV_ISA_Zbkx : boolean;
        RISCV_ISA_Zbs : boolean;
        RISCV_ISA_Zfinx : boolean;
        RISCV_ISA_Zicntr : boolean;
        RISCV_ISA_Zicond : boolean;
        RISCV_ISA_Zihpm : boolean;
        RISCV_ISA_Zkn : boolean;
        RISCV_ISA_Zknd : boolean;
        RISCV_ISA_Zkne : boolean;
        RISCV_ISA_Zknh : boolean;
        RISCV_ISA_Zks : boolean;
        RISCV_ISA_Zksed : boolean;
        RISCV_ISA_Zksh : boolean;
        RISCV_ISA_Zkt : boolean;
        RISCV_ISA_Zmmul : boolean;
        RISCV_ISA_Zxcfu : boolean;
        RISCV_ISA_Sdext : boolean;
        RISCV_ISA_Sdtrig : boolean;
        RISCV_ISA_Smpmp : boolean;
        CPU_FAST_MUL_EN : boolean;
        CPU_FAST_SHIFT_EN : boolean;
        CPU_RF_HW_RST_EN : boolean
    );
    port (
        clk_i : in std_ulogic;
        rstn_i : in std_ulogic;
        ctrl_o : out ctrl_bus_t;
        frontend_i : in if_bus_t;
        pmp_fault_i : in std_ulogic;
        alu_cp_done_i : in std_ulogic;
        alu_cmp_i : in std_ulogic_vector(1 downto 0);
        alu_add_i : in std_ulogic_vector(XLEN-1 downto 0);
        rf_rs1_i : in std_ulogic_vector(XLEN-1 downto 0);
        csr_rdata_o : out std_ulogic_vector(XLEN-1 downto 0);
        xcsr_rdata_i : in std_ulogic_vector(XLEN-1 downto 0);
        irq_dbg_i : in std_ulogic;
        irq_machine_i : in std_ulogic_vector(2 downto 0);
        irq_fast_i : in std_ulogic_vector(15 downto 0);
        lsu_wait_i : in std_ulogic;
        lsu_mar_i : in std_ulogic_vector(XLEN-1 downto 0);
        lsu_err_i : in std_ulogic_vector(3 downto 0);
        mem_sync_i : in std_ulogic
    );
end entity neorv32_cpu_control;